`timescale 1us / 1us
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/20/2024 04:19:42 PM
// Design Name: 
// Module Name: example_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module example_sim();
   
    reg clock_;
    always #5 clock_ = ~clock_;
    
    reg reset_;
    

    wire [31:0] cosout_;
    reg [31:0] x0_, y0_, z0_;
    wire [31:0] xn_, yn_, zn_;

    CORDIC cordicdut(
    .clock(clock_),
    .reset(reset_),
    .io_in_x0(x0_),
    .io_in_y0(y0_),
    .io_in_z0(z0_),
    .io_out_x(xn_),
    .io_out_y(yn_),
    .io_out_z(zn_)

    );
/*
Cos cosdut(
	.clock(clock_),
	.reset(reset_),
	.io_in(z0_),
	.io_out(cosout_));
*/


integer idx;
integer cyclecount;
 initial begin
    clock_ = 1'b0;
    reset_ = 1'b1;
	#10;


    reset_ = 1'b0;
    x0_ = 32'd1058764014;
	//x0_ = 32'h3f800000;
    y0_ = 32'h00000000;
    z0_ = 32'h3f490fdb;

#10;
z0_ = 32'hbfc90fdb; #10; //cos(-1.570796)=-0.000000, sin(-1.570796)=-1.000000
z0_ = 32'hbfc5eb9c; #10; //cos(-1.546253)=0.024541, sin(-1.546253)=-0.999699
z0_ = 32'hbfc2c75c; #10; //cos(-1.521709)=0.049068, sin(-1.521709)=-0.998795
z0_ = 32'hbfbfa31d; #10; //cos(-1.497165)=0.073564, sin(-1.497165)=-0.997290
z0_ = 32'hbfbc7edd; #10; //cos(-1.472622)=0.098017, sin(-1.472622)=-0.995185
z0_ = 32'hbfb95a9e; #10; //cos(-1.448078)=0.122411, sin(-1.448078)=-0.992480
z0_ = 32'hbfb6365e; #10; //cos(-1.423534)=0.146730, sin(-1.423534)=-0.989177
z0_ = 32'hbfb3121f; #10; //cos(-1.398991)=0.170962, sin(-1.398991)=-0.985278
z0_ = 32'hbfafede0; #10; //cos(-1.374447)=0.195090, sin(-1.374447)=-0.980785
z0_ = 32'hbfacc9a0; #10; //cos(-1.349903)=0.219101, sin(-1.349903)=-0.975702
z0_ = 32'hbfa9a561; #10; //cos(-1.325359)=0.242980, sin(-1.325359)=-0.970031
z0_ = 32'hbfa68121; #10; //cos(-1.300816)=0.266713, sin(-1.300816)=-0.963776
z0_ = 32'hbfa35ce2; #10; //cos(-1.276272)=0.290285, sin(-1.276272)=-0.956940
z0_ = 32'hbfa038a2; #10; //cos(-1.251728)=0.313682, sin(-1.251728)=-0.949528
z0_ = 32'hbf9d1463; #10; //cos(-1.227185)=0.336890, sin(-1.227185)=-0.941544
z0_ = 32'hbf99f024; #10; //cos(-1.202641)=0.359895, sin(-1.202641)=-0.932993
z0_ = 32'hbf96cbe4; #10; //cos(-1.178097)=0.382683, sin(-1.178097)=-0.923880
z0_ = 32'hbf93a7a5; #10; //cos(-1.153554)=0.405241, sin(-1.153554)=-0.914210
z0_ = 32'hbf908366; #10; //cos(-1.129010)=0.427555, sin(-1.129010)=-0.903989
z0_ = 32'hbf8d5f26; #10; //cos(-1.104466)=0.449611, sin(-1.104466)=-0.893224
z0_ = 32'hbf8a3ae6; #10; //cos(-1.079922)=0.471397, sin(-1.079922)=-0.881921
z0_ = 32'hbf8716a7; #10; //cos(-1.055379)=0.492898, sin(-1.055379)=-0.870087
z0_ = 32'hbf83f268; #10; //cos(-1.030835)=0.514103, sin(-1.030835)=-0.857729
z0_ = 32'hbf80ce28; #10; //cos(-1.006291)=0.534998, sin(-1.006291)=-0.844854
z0_ = 32'hbf7b53d2; #10; //cos(-0.981748)=0.555570, sin(-0.981748)=-0.831470
z0_ = 32'hbf750b53; #10; //cos(-0.957204)=0.575808, sin(-0.957204)=-0.817585
z0_ = 32'hbf6ec2d4; #10; //cos(-0.932660)=0.595699, sin(-0.932660)=-0.803208
z0_ = 32'hbf687a55; #10; //cos(-0.908117)=0.615232, sin(-0.908117)=-0.788346
z0_ = 32'hbf6231d6; #10; //cos(-0.883573)=0.634393, sin(-0.883573)=-0.773010
z0_ = 32'hbf5be958; #10; //cos(-0.859029)=0.653173, sin(-0.859029)=-0.757209
z0_ = 32'hbf55a0d9; #10; //cos(-0.834486)=0.671559, sin(-0.834486)=-0.740951
z0_ = 32'hbf4f585a; #10; //cos(-0.809942)=0.689541, sin(-0.809942)=-0.724247
z0_ = 32'hbf490fdb; #10; //cos(-0.785398)=0.707107, sin(-0.785398)=-0.707107
z0_ = 32'hbf42c75c; #10; //cos(-0.760854)=0.724247, sin(-0.760854)=-0.689541
z0_ = 32'hbf3c7edd; #10; //cos(-0.736311)=0.740951, sin(-0.736311)=-0.671559
z0_ = 32'hbf36365e; #10; //cos(-0.711767)=0.757209, sin(-0.711767)=-0.653173
z0_ = 32'hbf2fede0; #10; //cos(-0.687223)=0.773010, sin(-0.687223)=-0.634393
z0_ = 32'hbf29a561; #10; //cos(-0.662680)=0.788346, sin(-0.662680)=-0.615232
z0_ = 32'hbf235ce2; #10; //cos(-0.638136)=0.803208, sin(-0.638136)=-0.595699
z0_ = 32'hbf1d1463; #10; //cos(-0.613592)=0.817585, sin(-0.613592)=-0.575808
z0_ = 32'hbf16cbe4; #10; //cos(-0.589049)=0.831470, sin(-0.589049)=-0.555570
z0_ = 32'hbf108366; #10; //cos(-0.564505)=0.844854, sin(-0.564505)=-0.534998
z0_ = 32'hbf0a3ae6; #10; //cos(-0.539961)=0.857729, sin(-0.539961)=-0.514103
z0_ = 32'hbf03f268; #10; //cos(-0.515418)=0.870087, sin(-0.515418)=-0.492898
z0_ = 32'hbefb53d0; #10; //cos(-0.490874)=0.881921, sin(-0.490874)=-0.471397
z0_ = 32'hbeeec2d4; #10; //cos(-0.466330)=0.893224, sin(-0.466330)=-0.449611
z0_ = 32'hbee231d8; #10; //cos(-0.441787)=0.903989, sin(-0.441787)=-0.427555
z0_ = 32'hbed5a0d8; #10; //cos(-0.417243)=0.914210, sin(-0.417243)=-0.405241
z0_ = 32'hbec90fdc; #10; //cos(-0.392699)=0.923880, sin(-0.392699)=-0.382683
z0_ = 32'hbebc7edc; #10; //cos(-0.368155)=0.932993, sin(-0.368155)=-0.359895
z0_ = 32'hbeafede0; #10; //cos(-0.343612)=0.941544, sin(-0.343612)=-0.336890
z0_ = 32'hbea35ce0; #10; //cos(-0.319068)=0.949528, sin(-0.319068)=-0.313682
z0_ = 32'hbe96cbe4; #10; //cos(-0.294524)=0.956940, sin(-0.294524)=-0.290285
z0_ = 32'hbe8a3ae8; #10; //cos(-0.269981)=0.963776, sin(-0.269981)=-0.266713
z0_ = 32'hbe7b53d0; #10; //cos(-0.245437)=0.970031, sin(-0.245437)=-0.242980
z0_ = 32'hbe6231d8; #10; //cos(-0.220893)=0.975702, sin(-0.220893)=-0.219101
z0_ = 32'hbe490fd8; #10; //cos(-0.196350)=0.980785, sin(-0.196350)=-0.195090
z0_ = 32'hbe2fede0; #10; //cos(-0.171806)=0.985278, sin(-0.171806)=-0.170962
z0_ = 32'hbe16cbe8; #10; //cos(-0.147262)=0.989177, sin(-0.147262)=-0.146731
z0_ = 32'hbdfb53d0; #10; //cos(-0.122718)=0.992480, sin(-0.122718)=-0.122411
z0_ = 32'hbdc90fe0; #10; //cos(-0.098175)=0.995185, sin(-0.098175)=-0.098017
z0_ = 32'hbd96cbe0; #10; //cos(-0.073631)=0.997290, sin(-0.073631)=-0.073565
z0_ = 32'hbd490fe0; #10; //cos(-0.049087)=0.998795, sin(-0.049087)=-0.049068
z0_ = 32'hbcc90fc0; #10; //cos(-0.024544)=0.999699, sin(-0.024544)=-0.024541
z0_ = 32'h00000000; #10; //cos(0.000000)=1.000000, sin(0.000000)=0.000000
z0_ = 32'h3cc90fc0; #10; //cos(0.024544)=0.999699, sin(0.024544)=0.024541
z0_ = 32'h3d490fe0; #10; //cos(0.049087)=0.998795, sin(0.049087)=0.049068
z0_ = 32'h3d96cbe0; #10; //cos(0.073631)=0.997290, sin(0.073631)=0.073565
z0_ = 32'h3dc90fe0; #10; //cos(0.098175)=0.995185, sin(0.098175)=0.098017
z0_ = 32'h3dfb53d0; #10; //cos(0.122718)=0.992480, sin(0.122718)=0.122411
z0_ = 32'h3e16cbe8; #10; //cos(0.147262)=0.989177, sin(0.147262)=0.146731
z0_ = 32'h3e2fede0; #10; //cos(0.171806)=0.985278, sin(0.171806)=0.170962
z0_ = 32'h3e490fd8; #10; //cos(0.196350)=0.980785, sin(0.196350)=0.195090
z0_ = 32'h3e6231d8; #10; //cos(0.220893)=0.975702, sin(0.220893)=0.219101
z0_ = 32'h3e7b53d0; #10; //cos(0.245437)=0.970031, sin(0.245437)=0.242980
z0_ = 32'h3e8a3ae8; #10; //cos(0.269981)=0.963776, sin(0.269981)=0.266713
z0_ = 32'h3e96cbe4; #10; //cos(0.294524)=0.956940, sin(0.294524)=0.290285
z0_ = 32'h3ea35ce0; #10; //cos(0.319068)=0.949528, sin(0.319068)=0.313682
z0_ = 32'h3eafede0; #10; //cos(0.343612)=0.941544, sin(0.343612)=0.336890
z0_ = 32'h3ebc7edc; #10; //cos(0.368155)=0.932993, sin(0.368155)=0.359895
z0_ = 32'h3ec90fdc; #10; //cos(0.392699)=0.923880, sin(0.392699)=0.382683
z0_ = 32'h3ed5a0d8; #10; //cos(0.417243)=0.914210, sin(0.417243)=0.405241
z0_ = 32'h3ee231d4; #10; //cos(0.441786)=0.903989, sin(0.441786)=0.427555
z0_ = 32'h3eeec2d4; #10; //cos(0.466330)=0.893224, sin(0.466330)=0.449611
z0_ = 32'h3efb53d4; #10; //cos(0.490874)=0.881921, sin(0.490874)=0.471397
z0_ = 32'h3f03f266; #10; //cos(0.515417)=0.870087, sin(0.515417)=0.492898
z0_ = 32'h3f0a3ae6; #10; //cos(0.539961)=0.857729, sin(0.539961)=0.514103
z0_ = 32'h3f108366; #10; //cos(0.564505)=0.844854, sin(0.564505)=0.534998
z0_ = 32'h3f16cbe6; #10; //cos(0.589049)=0.831470, sin(0.589049)=0.555570
z0_ = 32'h3f1d1462; #10; //cos(0.613592)=0.817585, sin(0.613592)=0.575808
z0_ = 32'h3f235ce2; #10; //cos(0.638136)=0.803208, sin(0.638136)=0.595699
z0_ = 32'h3f29a562; #10; //cos(0.662680)=0.788346, sin(0.662680)=0.615232
z0_ = 32'h3f2fedde; #10; //cos(0.687223)=0.773010, sin(0.687223)=0.634393
z0_ = 32'h3f36365e; #10; //cos(0.711767)=0.757209, sin(0.711767)=0.653173
z0_ = 32'h3f3c7ede; #10; //cos(0.736311)=0.740951, sin(0.736311)=0.671559
z0_ = 32'h3f42c75e; #10; //cos(0.760855)=0.724247, sin(0.760855)=0.689541
z0_ = 32'h3f490fda; #10; //cos(0.785398)=0.707107, sin(0.785398)=0.707107
z0_ = 32'h3f4f585a; #10; //cos(0.809942)=0.689541, sin(0.809942)=0.724247
z0_ = 32'h3f55a0da; #10; //cos(0.834486)=0.671559, sin(0.834486)=0.740951
z0_ = 32'h3f5be956; #10; //cos(0.859029)=0.653173, sin(0.859029)=0.757209
z0_ = 32'h3f6231d6; #10; //cos(0.883573)=0.634393, sin(0.883573)=0.773010
z0_ = 32'h3f687a56; #10; //cos(0.908117)=0.615232, sin(0.908117)=0.788346
z0_ = 32'h3f6ec2d6; #10; //cos(0.932660)=0.595699, sin(0.932660)=0.803208
z0_ = 32'h3f750b52; #10; //cos(0.957204)=0.575808, sin(0.957204)=0.817585
z0_ = 32'h3f7b53d2; #10; //cos(0.981748)=0.555570, sin(0.981748)=0.831470
z0_ = 32'h3f80ce29; #10; //cos(1.006292)=0.534998, sin(1.006292)=0.844854
z0_ = 32'h3f83f267; #10; //cos(1.030835)=0.514103, sin(1.030835)=0.857729
z0_ = 32'h3f8716a7; #10; //cos(1.055379)=0.492898, sin(1.055379)=0.870087
z0_ = 32'h3f8a3ae7; #10; //cos(1.079923)=0.471397, sin(1.079923)=0.881921
z0_ = 32'h3f8d5f25; #10; //cos(1.104466)=0.449611, sin(1.104466)=0.893224
z0_ = 32'h3f908365; #10; //cos(1.129010)=0.427555, sin(1.129010)=0.903989
z0_ = 32'h3f93a7a5; #10; //cos(1.153554)=0.405241, sin(1.153554)=0.914210
z0_ = 32'h3f96cbe5; #10; //cos(1.178097)=0.382683, sin(1.178097)=0.923880
z0_ = 32'h3f99f023; #10; //cos(1.202641)=0.359895, sin(1.202641)=0.932993
z0_ = 32'h3f9d1463; #10; //cos(1.227185)=0.336890, sin(1.227185)=0.941544
z0_ = 32'h3fa038a3; #10; //cos(1.251728)=0.313682, sin(1.251728)=0.949528
z0_ = 32'h3fa35ce1; #10; //cos(1.276272)=0.290285, sin(1.276272)=0.956940
z0_ = 32'h3fa68121; #10; //cos(1.300816)=0.266713, sin(1.300816)=0.963776
z0_ = 32'h3fa9a561; #10; //cos(1.325359)=0.242980, sin(1.325359)=0.970031
z0_ = 32'h3facc9a1; #10; //cos(1.349903)=0.219101, sin(1.349903)=0.975702
z0_ = 32'h3fafeddf; #10; //cos(1.374447)=0.195090, sin(1.374447)=0.980785
z0_ = 32'h3fb3121f; #10; //cos(1.398991)=0.170962, sin(1.398991)=0.985278
z0_ = 32'h3fb6365f; #10; //cos(1.423534)=0.146730, sin(1.423534)=0.989177
z0_ = 32'h3fb95a9d; #10; //cos(1.448078)=0.122411, sin(1.448078)=0.992480
z0_ = 32'h3fbc7edd; #10; //cos(1.472622)=0.098017, sin(1.472622)=0.995185
z0_ = 32'h3fbfa31d; #10; //cos(1.497165)=0.073564, sin(1.497165)=0.997290
z0_ = 32'h3fc2c75d; #10; //cos(1.521709)=0.049068, sin(1.521709)=0.998795
z0_ = 32'h3fc5eb9b; #10; //cos(1.546253)=0.024541, sin(1.546253)=0.999699
z0_ = 32'h3fc90fdb; #10; //cos(1.570796)=-0.000000, sin(1.570796)=1.000000

    
 end
    
endmodule

