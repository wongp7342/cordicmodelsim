`timescale 1us / 1us

module example_sim();
    reg clock_;
    always #5 clock_ = ~clock_;
    reg reset_;
    

    wire [31:0] cosout_, sinout_;
    reg [31:0] x0_, y0_, z0_;

Sin sindut(
	.clock(clock_),
	.reset(reset_),
	.io_in(z0_),
	.io_out(sinout_));


integer idx;
integer cyclecount;
 initial begin

    clock_ = 1'b0;
    reset_ = 1'b1;
	#10;

    reset_ = 1'b0;
z0_ = 32'hc0c90fdb; #10; //cos(-6.283185)=1.000000, sin(-6.283185)=-0.000000
z0_ = 32'hc0c2c75c; #10; //cos(-6.086836)=0.980785, sin(-6.086836)=0.195090
z0_ = 32'hc0bc7edd; #10; //cos(-5.890486)=0.923880, sin(-5.890486)=0.382683
z0_ = 32'hc0b6365e; #10; //cos(-5.694137)=0.831470, sin(-5.694137)=0.555570
z0_ = 32'hc0afede0; #10; //cos(-5.497787)=0.707107, sin(-5.497787)=0.707107
z0_ = 32'hc0a9a561; #10; //cos(-5.301438)=0.555570, sin(-5.301438)=0.831469
z0_ = 32'hc0a35ce2; #10; //cos(-5.105088)=0.382684, sin(-5.105088)=0.923879
z0_ = 32'hc09d1463; #10; //cos(-4.908739)=0.195090, sin(-4.908739)=0.980785
z0_ = 32'hc096cbe4; #10; //cos(-4.712389)=0.000000, sin(-4.712389)=1.000000
z0_ = 32'hc0908366; #10; //cos(-4.516040)=-0.195090, sin(-4.516040)=0.980785
z0_ = 32'hc08a3ae6; #10; //cos(-4.319690)=-0.382684, sin(-4.319690)=0.923880
z0_ = 32'hc083f268; #10; //cos(-4.123341)=-0.555570, sin(-4.123341)=0.831470
z0_ = 32'hc07b53d2; #10; //cos(-3.926991)=-0.707107, sin(-3.926991)=0.707107
z0_ = 32'hc06ec2d4; #10; //cos(-3.730641)=-0.831470, sin(-3.730641)=0.555570
z0_ = 32'hc06231d6; #10; //cos(-3.534292)=-0.923880, sin(-3.534292)=0.382683
z0_ = 32'hc055a0d9; #10; //cos(-3.337942)=-0.980785, sin(-3.337942)=0.195090
z0_ = 32'hc0490fdb; #10; //cos(-3.141593)=-1.000000, sin(-3.141593)=0.000000
z0_ = 32'hc03c7edd; #10; //cos(-2.945243)=-0.980785, sin(-2.945243)=-0.195090
z0_ = 32'hc02fede0; #10; //cos(-2.748894)=-0.923880, sin(-2.748894)=-0.382683
z0_ = 32'hc0235ce2; #10; //cos(-2.552544)=-0.831470, sin(-2.552544)=-0.555570
z0_ = 32'hc016cbe4; #10; //cos(-2.356194)=-0.707107, sin(-2.356194)=-0.707107
z0_ = 32'hc00a3ae6; #10; //cos(-2.159845)=-0.555570, sin(-2.159845)=-0.831470
z0_ = 32'hbffb53d0; #10; //cos(-1.963495)=-0.382683, sin(-1.963495)=-0.923880
z0_ = 32'hbfe231d8; #10; //cos(-1.767146)=-0.195091, sin(-1.767146)=-0.980785
z0_ = 32'hbfc90fdc; #10; //cos(-1.570796)=-0.000000, sin(-1.570796)=-1.000000
z0_ = 32'hbfafede0; #10; //cos(-1.374447)=0.195090, sin(-1.374447)=-0.980785
z0_ = 32'hbf96cbe4; #10; //cos(-1.178097)=0.382683, sin(-1.178097)=-0.923880
z0_ = 32'hbf7b53d0; #10; //cos(-0.981748)=0.555570, sin(-0.981748)=-0.831470
z0_ = 32'hbf490fd8; #10; //cos(-0.785398)=0.707107, sin(-0.785398)=-0.707107
z0_ = 32'hbf16cbe8; #10; //cos(-0.589049)=0.831469, sin(-0.589049)=-0.555570
z0_ = 32'hbec90fe0; #10; //cos(-0.392699)=0.923879, sin(-0.392699)=-0.382684
z0_ = 32'hbe490fe0; #10; //cos(-0.196350)=0.980785, sin(-0.196350)=-0.195090
z0_ = 32'h00000000; #10; //cos(0.000000)=1.000000, sin(0.000000)=0.000000
z0_ = 32'h3e490fe0; #10; //cos(0.196350)=0.980785, sin(0.196350)=0.195090
z0_ = 32'h3ec90fe0; #10; //cos(0.392699)=0.923879, sin(0.392699)=0.382684
z0_ = 32'h3f16cbe8; #10; //cos(0.589049)=0.831469, sin(0.589049)=0.555570
z0_ = 32'h3f490fd8; #10; //cos(0.785398)=0.707107, sin(0.785398)=0.707107
z0_ = 32'h3f7b53d0; #10; //cos(0.981748)=0.555570, sin(0.981748)=0.831470
z0_ = 32'h3f96cbe4; #10; //cos(1.178097)=0.382683, sin(1.178097)=0.923880
z0_ = 32'h3fafede0; #10; //cos(1.374447)=0.195090, sin(1.374447)=0.980785
z0_ = 32'h3fc90fdc; #10; //cos(1.570796)=-0.000000, sin(1.570796)=1.000000
z0_ = 32'h3fe231d4; #10; //cos(1.767146)=-0.195090, sin(1.767146)=0.980785
z0_ = 32'h3ffb53d4; #10; //cos(1.963496)=-0.382684, sin(1.963496)=0.923879
z0_ = 32'h400a3ae6; #10; //cos(2.159845)=-0.555570, sin(2.159845)=0.831470
z0_ = 32'h4016cbe6; #10; //cos(2.356195)=-0.707107, sin(2.356195)=0.707106
z0_ = 32'h40235ce2; #10; //cos(2.552544)=-0.831470, sin(2.552544)=0.555570
z0_ = 32'h402fedde; #10; //cos(2.748893)=-0.923879, sin(2.748893)=0.382684
z0_ = 32'h403c7ede; #10; //cos(2.945243)=-0.980785, sin(2.945243)=0.195090
z0_ = 32'h40490fda; #10; //cos(3.141593)=-1.000000, sin(3.141593)=0.000000
z0_ = 32'h4055a0da; #10; //cos(3.337943)=-0.980785, sin(3.337943)=-0.195091
z0_ = 32'h406231d6; #10; //cos(3.534292)=-0.923880, sin(3.534292)=-0.382683
z0_ = 32'h406ec2d6; #10; //cos(3.730642)=-0.831469, sin(3.730642)=-0.555571
z0_ = 32'h407b53d2; #10; //cos(3.926991)=-0.707107, sin(3.926991)=-0.707107
z0_ = 32'h4083f267; #10; //cos(4.123340)=-0.555570, sin(4.123340)=-0.831469
z0_ = 32'h408a3ae7; #10; //cos(4.319690)=-0.382683, sin(4.319690)=-0.923880
z0_ = 32'h40908365; #10; //cos(4.516039)=-0.195090, sin(4.516039)=-0.980785
z0_ = 32'h4096cbe5; #10; //cos(4.712389)=0.000000, sin(4.712389)=-1.000000
z0_ = 32'h409d1463; #10; //cos(4.908739)=0.195090, sin(4.908739)=-0.980785
z0_ = 32'h40a35ce1; #10; //cos(5.105088)=0.382683, sin(5.105088)=-0.923880
z0_ = 32'h40a9a561; #10; //cos(5.301438)=0.555570, sin(5.301438)=-0.831469
z0_ = 32'h40afeddf; #10; //cos(5.497787)=0.707107, sin(5.497787)=-0.707107
z0_ = 32'h40b6365f; #10; //cos(5.694137)=0.831470, sin(5.694137)=-0.555570
z0_ = 32'h40bc7edd; #10; //cos(5.890486)=0.923880, sin(5.890486)=-0.382683
z0_ = 32'h40c2c75d; #10; //cos(6.086836)=0.980785, sin(6.086836)=-0.195090
z0_ = 32'h40c90fdb; #10; //cos(6.283185)=1.000000, sin(6.283185)=0.000000

    
 end
    
endmodule

