`timescale 1us / 1us

module example_sim();
	reg [31:0] clockcount_;
    reg clock_;
    always #5 clock_ = ~clock_;
    reg reset_;
    always #10 clockcount_ = clockcount_ + 1;

    wire [31:0] cosout_, sinout_;
    reg [31:0] x0_, y0_, z0_;

Sin sindut(
	.clock(clock_),
	.reset(reset_),
	.io_in(z0_),
	.io_out(sinout_));


integer idx;
integer cyclecount;
initial begin
	clockcount_ = 32'd0;
    clock_ = 1'b1;
    reset_ = 1'b1;
	#10;

    reset_ = 1'b0;
    #10;
    /* Though they look like common angles in degrees, the angles in 
		the comments are in fact radians, NOT degrees
    */
    z0_ = 32'hc27b53d2; #10; //cos(-62.831856)=1.000000, sin(-62.831856)=-0.000003
	z0_ = 32'hc2737933; #10; //cos(-60.868359)=-0.382683, sin(-60.868359)=0.923880
	z0_ = 32'hc26b9e94; #10; //cos(-58.904861)=-0.707106, sin(-58.904861)=-0.707107
	z0_ = 32'hc263c3f6; #10; //cos(-56.941368)=0.923879, sin(-56.941368)=-0.382685
	z0_ = 32'hc25be958; #10; //cos(-54.977875)=0.000003, sin(-54.977875)=1.000000
	z0_ = 32'hc2540eb9; #10; //cos(-53.014378)=-0.923880, sin(-53.014378)=-0.382682
	z0_ = 32'hc24c341a; #10; //cos(-51.050880)=0.707107, sin(-51.050880)=-0.707107
	z0_ = 32'hc244597c; #10; //cos(-49.087387)=0.382685, sin(-49.087387)=0.923879
	z0_ = 32'hc23c7edd; #10; //cos(-47.123890)=-1.000000, sin(-47.123890)=0.000000
	z0_ = 32'hc234a440; #10; //cos(-45.160400)=0.382678, sin(-45.160400)=-0.923882
	z0_ = 32'hc22cc9a0; #10; //cos(-43.196899)=0.707107, sin(-43.196899)=0.707106
	z0_ = 32'hc224ef02; #10; //cos(-41.233406)=-0.923879, sin(-41.233406)=0.382686
	z0_ = 32'hc21d1463; #10; //cos(-39.269909)=-0.000001, sin(-39.269909)=-1.000000
	z0_ = 32'hc21539c4; #10; //cos(-37.306412)=0.923879, sin(-37.306412)=0.382684
	z0_ = 32'hc20d5f26; #10; //cos(-35.342918)=-0.707106, sin(-35.342918)=0.707108
	z0_ = 32'hc2058488; #10; //cos(-33.379425)=-0.382686, sin(-33.379425)=-0.923878
	z0_ = 32'hc1fb53d2; #10; //cos(-31.415928)=1.000000, sin(-31.415928)=-0.000001
	z0_ = 32'hc1eb9e94; #10; //cos(-29.452431)=-0.382684, sin(-29.452431)=0.923879
	z0_ = 32'hc1dbe958; #10; //cos(-27.488937)=-0.707108, sin(-27.488937)=-0.707106
	z0_ = 32'hc1cc341a; #10; //cos(-25.525440)=0.923880, sin(-25.525440)=-0.382683
	z0_ = 32'hc1bc7edd; #10; //cos(-23.561945)=0.000000, sin(-23.561945)=1.000000
	z0_ = 32'hc1acc9a0; #10; //cos(-21.598450)=-0.923880, sin(-21.598450)=-0.382683
	z0_ = 32'hc19d1462; #10; //cos(-19.634953)=0.707108, sin(-19.634953)=-0.707106
	z0_ = 32'hc18d5f27; #10; //cos(-17.671461)=0.382686, sin(-17.671461)=0.923879
	z0_ = 32'hc17b53d3; #10; //cos(-15.707965)=-1.000000, sin(-15.707965)=0.000002
	z0_ = 32'hc15be958; #10; //cos(-13.744469)=0.382683, sin(-13.744469)=-0.923880
	z0_ = 32'hc13c7edd; #10; //cos(-11.780972)=0.707107, sin(-11.780972)=0.707107
	z0_ = 32'hc11d1462; #10; //cos(-9.817476)=-0.923880, sin(-9.817476)=0.382683
	z0_ = 32'hc0fb53ce; #10; //cos(-7.853980)=0.000002, sin(-7.853980)=-1.000000
	z0_ = 32'hc0bc7ee2; #10; //cos(-5.890489)=0.923880, sin(-5.890489)=0.382681
	z0_ = 32'hc07b53d8; #10; //cos(-3.926992)=-0.707106, sin(-3.926992)=0.707108
	z0_ = 32'hbffb53d8; #10; //cos(-1.963496)=-0.382684, sin(-1.963496)=-0.923879
	z0_ = 32'h00000000; #10; //cos(0.000000)=1.000000, sin(0.000000)=0.000000
	z0_ = 32'h3ffb53d8; #10; //cos(1.963496)=-0.382684, sin(1.963496)=0.923879
	z0_ = 32'h407b53d8; #10; //cos(3.926992)=-0.707106, sin(3.926992)=-0.707108
	z0_ = 32'h40bc7ee2; #10; //cos(5.890489)=0.923880, sin(5.890489)=-0.382681
	z0_ = 32'h40fb53ce; #10; //cos(7.853980)=0.000002, sin(7.853980)=1.000000
	z0_ = 32'h411d1462; #10; //cos(9.817476)=-0.923880, sin(9.817476)=-0.382683
	z0_ = 32'h413c7edd; #10; //cos(11.780972)=0.707107, sin(11.780972)=-0.707107
	z0_ = 32'h415be958; #10; //cos(13.744469)=0.382683, sin(13.744469)=0.923880
	z0_ = 32'h417b53d3; #10; //cos(15.707965)=-1.000000, sin(15.707965)=-0.000002
	z0_ = 32'h418d5f24; #10; //cos(17.671455)=0.382680, sin(17.671455)=-0.923881
	z0_ = 32'h419d1464; #10; //cos(19.634956)=0.707105, sin(19.634956)=0.707108
	z0_ = 32'h41acc9a0; #10; //cos(21.598450)=-0.923880, sin(21.598450)=0.382683
	z0_ = 32'h41bc7ee0; #10; //cos(23.561951)=0.000006, sin(23.561951)=-1.000000
	z0_ = 32'h41cc341a; #10; //cos(25.525440)=0.923880, sin(25.525440)=0.382683
	z0_ = 32'h41dbe956; #10; //cos(27.488934)=-0.707105, sin(27.488934)=0.707108
	z0_ = 32'h41eb9e96; #10; //cos(29.452435)=-0.382680, sin(29.452435)=-0.923881
	z0_ = 32'h41fb53d0; #10; //cos(31.415924)=1.000000, sin(31.415924)=-0.000002
	z0_ = 32'h42058488; #10; //cos(33.379425)=-0.382686, sin(33.379425)=0.923878
	z0_ = 32'h420d5f26; #10; //cos(35.342918)=-0.707106, sin(35.342918)=-0.707108
	z0_ = 32'h421539c6; #10; //cos(37.306419)=0.923882, sin(37.306419)=-0.382677
	z0_ = 32'h421d1463; #10; //cos(39.269909)=-0.000001, sin(39.269909)=1.000000
	z0_ = 32'h4224ef01; #10; //cos(41.233402)=-0.923880, sin(41.233402)=-0.382682
	z0_ = 32'h422cc9a1; #10; //cos(43.196903)=0.707110, sin(43.196903)=-0.707104
	z0_ = 32'h4234a43e; #10; //cos(45.160393)=0.382685, sin(45.160393)=0.923879
	z0_ = 32'h423c7ede; #10; //cos(47.123894)=-1.000000, sin(47.123894)=-0.000004
	z0_ = 32'h4244597c; #10; //cos(49.087387)=0.382685, sin(49.087387)=-0.923879
	z0_ = 32'h424c3419; #10; //cos(51.050877)=0.707110, sin(51.050877)=0.707104
	z0_ = 32'h42540eb9; #10; //cos(53.014378)=-0.923880, sin(53.014378)=0.382682
	z0_ = 32'h425be957; #10; //cos(54.977871)=-0.000000, sin(54.977871)=-1.000000
	z0_ = 32'h4263c3f7; #10; //cos(56.941372)=0.923878, sin(56.941372)=0.382688
	z0_ = 32'h426b9e94; #10; //cos(58.904861)=-0.707106, sin(58.904861)=0.707107
	z0_ = 32'h42737934; #10; //cos(60.868362)=-0.382679, sin(60.868362)=-0.923881
	z0_ = 32'h427b53d2; #10; //cos(62.831856)=1.000000, sin(62.831856)=0.000003


    
end
    
endmodule

