module FloatToFixed32(
  input  [31:0] io_in,
  output [31:0] io_out
);
  wire [31:0] frac = {9'h0,io_in[22:0]}; // @[FixedPoint.scala 17:42]
  wire [7:0] exp = io_in[30:23]; // @[FixedPoint.scala 18:25]
  wire  sign = io_in[31]; // @[FixedPoint.scala 19:26]
  wire [7:0] shiftamt = exp - 8'h7f; // @[FixedPoint.scala 20:37]
  wire [31:0] _data_T_3 = frac | 32'h800000; // @[FixedPoint.scala 23:18]
  wire [36:0] _GEN_0 = {_data_T_3, 5'h0}; // @[FixedPoint.scala 23:40]
  wire [38:0] _data_T_4 = {{2'd0}, _GEN_0}; // @[FixedPoint.scala 23:40]
  wire [7:0] _data_T_8 = 8'sh0 - $signed(shiftamt); // @[FixedPoint.scala 23:63]
  wire [38:0] _data_T_9 = _data_T_4 >> _data_T_8; // @[FixedPoint.scala 23:48]
  wire [7:0] _data_T_13 = exp - 8'h7f; // @[FixedPoint.scala 24:62]
  wire [293:0] _GEN_1 = {{255'd0}, _data_T_4}; // @[FixedPoint.scala 24:48]
  wire [293:0] _data_T_14 = _GEN_1 << _data_T_13; // @[FixedPoint.scala 24:48]
  wire [293:0] data = shiftamt[7] ? {{255'd0}, _data_T_9} : _data_T_14; // @[FixedPoint.scala 22:17]
  wire [293:0] _io_out_T_3 = 294'h0 - data; // @[FixedPoint.scala 25:40]
  wire [293:0] _io_out_T_4 = sign ? _io_out_T_3 : data; // @[FixedPoint.scala 25:16]
  assign io_out = _io_out_T_4[31:0]; // @[FixedPoint.scala 25:10]
endmodule
module CLZ32(
  input  [31:0] io_in,
  output [4:0]  io_out
);
  wire [31:0] _bx_T = io_in & 32'hffff0000; // @[FixedPoint.scala 36:20]
  wire  _bx_T_1 = _bx_T == 32'h0; // @[FixedPoint.scala 36:37]
  wire [47:0] _bx_T_2 = {io_in, 16'h0}; // @[FixedPoint.scala 36:49]
  wire [47:0] bx = _bx_T == 32'h0 ? _bx_T_2 : {{16'd0}, io_in}; // @[FixedPoint.scala 36:15]
  wire [47:0] _cx_T = bx & 48'hff000000; // @[FixedPoint.scala 37:20]
  wire  _cx_T_1 = _cx_T == 48'h0; // @[FixedPoint.scala 37:37]
  wire [55:0] _cx_T_2 = {bx, 8'h0}; // @[FixedPoint.scala 37:49]
  wire [55:0] cx = _cx_T == 48'h0 ? _cx_T_2 : {{8'd0}, bx}; // @[FixedPoint.scala 37:15]
  wire [55:0] _dx_T = cx & 56'hf0000000; // @[FixedPoint.scala 38:20]
  wire  _dx_T_1 = _dx_T == 56'h0; // @[FixedPoint.scala 38:37]
  wire [59:0] _dx_T_2 = {cx, 4'h0}; // @[FixedPoint.scala 38:49]
  wire [59:0] dx = _dx_T == 56'h0 ? _dx_T_2 : {{4'd0}, cx}; // @[FixedPoint.scala 38:15]
  wire [59:0] _ex_T = dx & 60'hc0000000; // @[FixedPoint.scala 39:20]
  wire  _ex_T_1 = _ex_T == 60'h0; // @[FixedPoint.scala 39:37]
  wire [61:0] _ex_T_2 = {dx, 2'h0}; // @[FixedPoint.scala 39:49]
  wire [61:0] ex = _ex_T == 60'h0 ? _ex_T_2 : {{2'd0}, dx}; // @[FixedPoint.scala 39:15]
  wire [3:0] _io_out_T_10 = {_bx_T_1,_cx_T_1,_dx_T_1,_ex_T_1}; // @[FixedPoint.scala 41:112]
  wire [61:0] _io_out_T_11 = ex & 62'h80000000; // @[FixedPoint.scala 42:44]
  assign io_out = {_io_out_T_10,_io_out_T_11 == 62'h0}; // @[FixedPoint.scala 42:36]
endmodule
module FixedToFloat32(
  input  [31:0] io_in,
  output [31:0] io_out
);
  wire [31:0] clz32_io_in; // @[FixedPoint.scala 62:21]
  wire [4:0] clz32_io_out; // @[FixedPoint.scala 62:21]
  wire [31:0] _data_T_2 = ~io_in; // @[FixedPoint.scala 59:35]
  wire [31:0] _data_T_4 = _data_T_2 + 32'h1; // @[FixedPoint.scala 59:50]
  wire [4:0] _leadingzeros_T = clz32_io_out; // @[FixedPoint.scala 65:47]
  wire [18:0] leadingzeros = {14'h0,_leadingzeros_T}; // @[FixedPoint.scala 65:32]
  wire [3:0] _exp_T_2 = 4'sh4 - 4'sh1; // @[FixedPoint.scala 67:16]
  wire [18:0] _exp_T_3 = {14'h0,_leadingzeros_T}; // @[FixedPoint.scala 67:38]
  wire [18:0] _GEN_0 = {{15{_exp_T_2[3]}},_exp_T_2}; // @[FixedPoint.scala 67:23]
  wire [18:0] _exp_T_6 = $signed(_GEN_0) - $signed(_exp_T_3); // @[FixedPoint.scala 67:23]
  wire [18:0] _exp_T_9 = $signed(_exp_T_6) + 19'sh7f; // @[FixedPoint.scala 67:46]
  wire [31:0] _frac_T = io_in[31] ? _data_T_4 : io_in; // @[FixedPoint.scala 68:19]
  wire [18:0] _frac_T_2 = leadingzeros + 19'h1; // @[FixedPoint.scala 68:43]
  wire [524318:0] _GEN_3 = {{524287{_frac_T[31]}},_frac_T}; // @[FixedPoint.scala 68:26]
  wire [524318:0] _frac_T_3 = $signed(_GEN_3) << _frac_T_2; // @[FixedPoint.scala 68:26]
  wire [5:0] _frac_T_5 = 6'h20 - 6'h17; // @[FixedPoint.scala 68:75]
  wire [524318:0] _frac_T_6 = $signed(_frac_T_3) >>> _frac_T_5; // @[FixedPoint.scala 68:66]
  wire [7:0] _io_out_T_1 = _exp_T_9[7:0]; // @[FixedPoint.scala 70:30]
  wire [8:0] _io_out_T_2 = {io_in[31],_io_out_T_1}; // @[FixedPoint.scala 70:23]
  wire [22:0] _io_out_T_3 = _frac_T_6[22:0]; // @[FixedPoint.scala 70:44]
  CLZ32 clz32 ( // @[FixedPoint.scala 62:21]
    .io_in(clz32_io_in),
    .io_out(clz32_io_out)
  );
  assign io_out = {_io_out_T_2,_io_out_T_3}; // @[FixedPoint.scala 70:37]
  assign clz32_io_in = io_in[31] ? _data_T_4 : io_in; // @[FixedPoint.scala 59:14]
endmodule
module CORDIC(
  input  [31:0] io_in_z0,
  input  [31:0] io_in_mode,
  output [31:0] io_out_x,
  output [1:0]  io_out_mode
);
  wire [31:0] tofixedx0_io_in; // @[CORDIC.scala 63:25]
  wire [31:0] tofixedx0_io_out; // @[CORDIC.scala 63:25]
  wire [31:0] tofixedy0_io_in; // @[CORDIC.scala 64:25]
  wire [31:0] tofixedy0_io_out; // @[CORDIC.scala 64:25]
  wire [31:0] tofloatxout_io_in; // @[CORDIC.scala 123:27]
  wire [31:0] tofloatxout_io_out; // @[CORDIC.scala 123:27]
  wire [31:0] tofloatyout_io_in; // @[CORDIC.scala 124:27]
  wire [31:0] tofloatyout_io_out; // @[CORDIC.scala 124:27]
  wire [31:0] tofloatzout_io_in; // @[CORDIC.scala 125:27]
  wire [31:0] tofloatzout_io_out; // @[CORDIC.scala 125:27]
  wire  _fxxterm_T = 32'sh0 > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_3 = 32'sh0 - $signed(tofixedx0_io_out); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm = 32'sh0 > $signed(io_in_z0) ? $signed(_fxxterm_T_3) : $signed(tofixedx0_io_out); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_3 = 32'sh0 - $signed(tofixedy0_io_out); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm = _fxxterm_T ? $signed(_fxyterm_T_3) : $signed(tofixedy0_io_out); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_2 = 32'h0 - 32'hc90fdb0; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_1_T = _fxxterm_T ? _fxthetaterm_T_2 : 32'hc90fdb0; // @[CORDIC.scala 116:44]
  wire [32:0] _theta_1_T_1 = {{1{_theta_1_T[31]}},_theta_1_T}; // @[CORDIC.scala 116:30]
  wire [31:0] theta_1 = _theta_1_T_1[31:0]; // @[CORDIC.scala 116:30]
  wire [31:0] x_1 = $signed(tofixedx0_io_out) - $signed(fxyterm); // @[CORDIC.scala 117:22]
  wire [31:0] y_1 = $signed(fxxterm) + $signed(tofixedy0_io_out); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_4 = $signed(theta_1) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_7 = 32'sh0 - $signed(x_1); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_1 = $signed(theta_1) > $signed(io_in_z0) ? $signed(_fxxterm_T_7) : $signed(x_1); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_7 = 32'sh0 - $signed(y_1); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_1 = _fxxterm_T_4 ? $signed(_fxyterm_T_7) : $signed(y_1); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_5 = 32'h0 - 32'h76b19c0; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_2_T = _fxxterm_T_4 ? _fxthetaterm_T_5 : 32'h76b19c0; // @[CORDIC.scala 116:44]
  wire [31:0] theta_2 = $signed(theta_1) + $signed(_theta_2_T); // @[CORDIC.scala 116:30]
  wire [30:0] _GEN_0 = fxyterm_1[31:1]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_2_T = {{1{_GEN_0[30]}},_GEN_0}; // @[CORDIC.scala 117:33]
  wire [31:0] x_2 = $signed(x_1) - $signed(_x_2_T); // @[CORDIC.scala 117:22]
  wire [30:0] _GEN_1 = fxxterm_1[31:1]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_2_T = {{1{_GEN_1[30]}},_GEN_1}; // @[CORDIC.scala 118:26]
  wire [31:0] y_2 = $signed(_y_2_T) + $signed(y_1); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_8 = $signed(theta_2) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_11 = 32'sh0 - $signed(x_2); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_2 = $signed(theta_2) > $signed(io_in_z0) ? $signed(_fxxterm_T_11) : $signed(x_2); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_11 = 32'sh0 - $signed(y_2); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_2 = _fxxterm_T_8 ? $signed(_fxyterm_T_11) : $signed(y_2); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_8 = 32'h0 - 32'h3eb6ec0; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_3_T = _fxxterm_T_8 ? _fxthetaterm_T_8 : 32'h3eb6ec0; // @[CORDIC.scala 116:44]
  wire [31:0] theta_3 = $signed(theta_2) + $signed(_theta_3_T); // @[CORDIC.scala 116:30]
  wire [29:0] _GEN_2 = fxyterm_2[31:2]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_3_T = {{2{_GEN_2[29]}},_GEN_2}; // @[CORDIC.scala 117:33]
  wire [31:0] x_3 = $signed(x_2) - $signed(_x_3_T); // @[CORDIC.scala 117:22]
  wire [29:0] _GEN_3 = fxxterm_2[31:2]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_3_T = {{2{_GEN_3[29]}},_GEN_3}; // @[CORDIC.scala 118:26]
  wire [31:0] y_3 = $signed(_y_3_T) + $signed(y_2); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_12 = $signed(theta_3) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_15 = 32'sh0 - $signed(x_3); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_3 = $signed(theta_3) > $signed(io_in_z0) ? $signed(_fxxterm_T_15) : $signed(x_3); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_15 = 32'sh0 - $signed(y_3); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_3 = _fxxterm_T_12 ? $signed(_fxyterm_T_15) : $signed(y_3); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_11 = 32'h0 - 32'h1fd5baa; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_4_T = _fxxterm_T_12 ? _fxthetaterm_T_11 : 32'h1fd5baa; // @[CORDIC.scala 116:44]
  wire [31:0] theta_4 = $signed(theta_3) + $signed(_theta_4_T); // @[CORDIC.scala 116:30]
  wire [28:0] _GEN_4 = fxyterm_3[31:3]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_4_T = {{3{_GEN_4[28]}},_GEN_4}; // @[CORDIC.scala 117:33]
  wire [31:0] x_4 = $signed(x_3) - $signed(_x_4_T); // @[CORDIC.scala 117:22]
  wire [28:0] _GEN_5 = fxxterm_3[31:3]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_4_T = {{3{_GEN_5[28]}},_GEN_5}; // @[CORDIC.scala 118:26]
  wire [31:0] y_4 = $signed(_y_4_T) + $signed(y_3); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_16 = $signed(theta_4) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_19 = 32'sh0 - $signed(x_4); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_4 = $signed(theta_4) > $signed(io_in_z0) ? $signed(_fxxterm_T_19) : $signed(x_4); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_19 = 32'sh0 - $signed(y_4); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_4 = _fxxterm_T_16 ? $signed(_fxyterm_T_19) : $signed(y_4); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_14 = 32'h0 - 32'hffaade; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_5_T = _fxxterm_T_16 ? _fxthetaterm_T_14 : 32'hffaade; // @[CORDIC.scala 116:44]
  wire [31:0] theta_5 = $signed(theta_4) + $signed(_theta_5_T); // @[CORDIC.scala 116:30]
  wire [27:0] _GEN_6 = fxyterm_4[31:4]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_5_T = {{4{_GEN_6[27]}},_GEN_6}; // @[CORDIC.scala 117:33]
  wire [31:0] x_5 = $signed(x_4) - $signed(_x_5_T); // @[CORDIC.scala 117:22]
  wire [27:0] _GEN_7 = fxxterm_4[31:4]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_5_T = {{4{_GEN_7[27]}},_GEN_7}; // @[CORDIC.scala 118:26]
  wire [31:0] y_5 = $signed(_y_5_T) + $signed(y_4); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_20 = $signed(theta_5) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_23 = 32'sh0 - $signed(x_5); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_5 = $signed(theta_5) > $signed(io_in_z0) ? $signed(_fxxterm_T_23) : $signed(x_5); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_23 = 32'sh0 - $signed(y_5); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_5 = _fxxterm_T_20 ? $signed(_fxyterm_T_23) : $signed(y_5); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_17 = 32'h0 - 32'h7ff557; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_6_T = _fxxterm_T_20 ? _fxthetaterm_T_17 : 32'h7ff557; // @[CORDIC.scala 116:44]
  wire [31:0] theta_6 = $signed(theta_5) + $signed(_theta_6_T); // @[CORDIC.scala 116:30]
  wire [26:0] _GEN_8 = fxyterm_5[31:5]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_6_T = {{5{_GEN_8[26]}},_GEN_8}; // @[CORDIC.scala 117:33]
  wire [31:0] x_6 = $signed(x_5) - $signed(_x_6_T); // @[CORDIC.scala 117:22]
  wire [26:0] _GEN_9 = fxxterm_5[31:5]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_6_T = {{5{_GEN_9[26]}},_GEN_9}; // @[CORDIC.scala 118:26]
  wire [31:0] y_6 = $signed(_y_6_T) + $signed(y_5); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_24 = $signed(theta_6) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_27 = 32'sh0 - $signed(x_6); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_6 = $signed(theta_6) > $signed(io_in_z0) ? $signed(_fxxterm_T_27) : $signed(x_6); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_27 = 32'sh0 - $signed(y_6); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_6 = _fxxterm_T_24 ? $signed(_fxyterm_T_27) : $signed(y_6); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_20 = 32'h0 - 32'h3ffeaa; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_7_T = _fxxterm_T_24 ? _fxthetaterm_T_20 : 32'h3ffeaa; // @[CORDIC.scala 116:44]
  wire [31:0] theta_7 = $signed(theta_6) + $signed(_theta_7_T); // @[CORDIC.scala 116:30]
  wire [25:0] _GEN_10 = fxyterm_6[31:6]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_7_T = {{6{_GEN_10[25]}},_GEN_10}; // @[CORDIC.scala 117:33]
  wire [31:0] x_7 = $signed(x_6) - $signed(_x_7_T); // @[CORDIC.scala 117:22]
  wire [25:0] _GEN_11 = fxxterm_6[31:6]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_7_T = {{6{_GEN_11[25]}},_GEN_11}; // @[CORDIC.scala 118:26]
  wire [31:0] y_7 = $signed(_y_7_T) + $signed(y_6); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_28 = $signed(theta_7) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_31 = 32'sh0 - $signed(x_7); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_7 = $signed(theta_7) > $signed(io_in_z0) ? $signed(_fxxterm_T_31) : $signed(x_7); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_31 = 32'sh0 - $signed(y_7); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_7 = _fxxterm_T_28 ? $signed(_fxyterm_T_31) : $signed(y_7); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_23 = 32'h0 - 32'h1fffd5; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_8_T = _fxxterm_T_28 ? _fxthetaterm_T_23 : 32'h1fffd5; // @[CORDIC.scala 116:44]
  wire [31:0] theta_8 = $signed(theta_7) + $signed(_theta_8_T); // @[CORDIC.scala 116:30]
  wire [24:0] _GEN_12 = fxyterm_7[31:7]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_8_T = {{7{_GEN_12[24]}},_GEN_12}; // @[CORDIC.scala 117:33]
  wire [31:0] x_8 = $signed(x_7) - $signed(_x_8_T); // @[CORDIC.scala 117:22]
  wire [24:0] _GEN_13 = fxxterm_7[31:7]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_8_T = {{7{_GEN_13[24]}},_GEN_13}; // @[CORDIC.scala 118:26]
  wire [31:0] y_8 = $signed(_y_8_T) + $signed(y_7); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_32 = $signed(theta_8) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_35 = 32'sh0 - $signed(x_8); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_8 = $signed(theta_8) > $signed(io_in_z0) ? $signed(_fxxterm_T_35) : $signed(x_8); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_35 = 32'sh0 - $signed(y_8); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_8 = _fxxterm_T_32 ? $signed(_fxyterm_T_35) : $signed(y_8); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_26 = 32'h0 - 32'hffffa; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_9_T = _fxxterm_T_32 ? _fxthetaterm_T_26 : 32'hffffa; // @[CORDIC.scala 116:44]
  wire [31:0] theta_9 = $signed(theta_8) + $signed(_theta_9_T); // @[CORDIC.scala 116:30]
  wire [23:0] _GEN_14 = fxyterm_8[31:8]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_9_T = {{8{_GEN_14[23]}},_GEN_14}; // @[CORDIC.scala 117:33]
  wire [31:0] x_9 = $signed(x_8) - $signed(_x_9_T); // @[CORDIC.scala 117:22]
  wire [23:0] _GEN_15 = fxxterm_8[31:8]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_9_T = {{8{_GEN_15[23]}},_GEN_15}; // @[CORDIC.scala 118:26]
  wire [31:0] y_9 = $signed(_y_9_T) + $signed(y_8); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_36 = $signed(theta_9) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_39 = 32'sh0 - $signed(x_9); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_9 = $signed(theta_9) > $signed(io_in_z0) ? $signed(_fxxterm_T_39) : $signed(x_9); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_39 = 32'sh0 - $signed(y_9); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_9 = _fxxterm_T_36 ? $signed(_fxyterm_T_39) : $signed(y_9); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_29 = 32'h0 - 32'h7ffff; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_10_T = _fxxterm_T_36 ? _fxthetaterm_T_29 : 32'h7ffff; // @[CORDIC.scala 116:44]
  wire [31:0] theta_10 = $signed(theta_9) + $signed(_theta_10_T); // @[CORDIC.scala 116:30]
  wire [22:0] _GEN_16 = fxyterm_9[31:9]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_10_T = {{9{_GEN_16[22]}},_GEN_16}; // @[CORDIC.scala 117:33]
  wire [31:0] x_10 = $signed(x_9) - $signed(_x_10_T); // @[CORDIC.scala 117:22]
  wire [22:0] _GEN_17 = fxxterm_9[31:9]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_10_T = {{9{_GEN_17[22]}},_GEN_17}; // @[CORDIC.scala 118:26]
  wire [31:0] y_10 = $signed(_y_10_T) + $signed(y_9); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_40 = $signed(theta_10) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_43 = 32'sh0 - $signed(x_10); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_10 = $signed(theta_10) > $signed(io_in_z0) ? $signed(_fxxterm_T_43) : $signed(x_10); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_43 = 32'sh0 - $signed(y_10); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_10 = _fxxterm_T_40 ? $signed(_fxyterm_T_43) : $signed(y_10); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_32 = 32'h0 - 32'h3ffff; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_11_T = _fxxterm_T_40 ? _fxthetaterm_T_32 : 32'h3ffff; // @[CORDIC.scala 116:44]
  wire [31:0] theta_11 = $signed(theta_10) + $signed(_theta_11_T); // @[CORDIC.scala 116:30]
  wire [21:0] _GEN_18 = fxyterm_10[31:10]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_11_T = {{10{_GEN_18[21]}},_GEN_18}; // @[CORDIC.scala 117:33]
  wire [31:0] x_11 = $signed(x_10) - $signed(_x_11_T); // @[CORDIC.scala 117:22]
  wire [21:0] _GEN_19 = fxxterm_10[31:10]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_11_T = {{10{_GEN_19[21]}},_GEN_19}; // @[CORDIC.scala 118:26]
  wire [31:0] y_11 = $signed(_y_11_T) + $signed(y_10); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_44 = $signed(theta_11) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_47 = 32'sh0 - $signed(x_11); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_11 = $signed(theta_11) > $signed(io_in_z0) ? $signed(_fxxterm_T_47) : $signed(x_11); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_47 = 32'sh0 - $signed(y_11); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_11 = _fxxterm_T_44 ? $signed(_fxyterm_T_47) : $signed(y_11); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_35 = 32'h0 - 32'h1ffff; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_12_T = _fxxterm_T_44 ? _fxthetaterm_T_35 : 32'h1ffff; // @[CORDIC.scala 116:44]
  wire [31:0] theta_12 = $signed(theta_11) + $signed(_theta_12_T); // @[CORDIC.scala 116:30]
  wire [20:0] _GEN_20 = fxyterm_11[31:11]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_12_T = {{11{_GEN_20[20]}},_GEN_20}; // @[CORDIC.scala 117:33]
  wire [31:0] x_12 = $signed(x_11) - $signed(_x_12_T); // @[CORDIC.scala 117:22]
  wire [20:0] _GEN_21 = fxxterm_11[31:11]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_12_T = {{11{_GEN_21[20]}},_GEN_21}; // @[CORDIC.scala 118:26]
  wire [31:0] y_12 = $signed(_y_12_T) + $signed(y_11); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_48 = $signed(theta_12) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_51 = 32'sh0 - $signed(x_12); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_12 = $signed(theta_12) > $signed(io_in_z0) ? $signed(_fxxterm_T_51) : $signed(x_12); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_51 = 32'sh0 - $signed(y_12); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_12 = _fxxterm_T_48 ? $signed(_fxyterm_T_51) : $signed(y_12); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_38 = 32'h0 - 32'h10000; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_13_T = _fxxterm_T_48 ? _fxthetaterm_T_38 : 32'h10000; // @[CORDIC.scala 116:44]
  wire [31:0] theta_13 = $signed(theta_12) + $signed(_theta_13_T); // @[CORDIC.scala 116:30]
  wire [19:0] _GEN_22 = fxyterm_12[31:12]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_13_T = {{12{_GEN_22[19]}},_GEN_22}; // @[CORDIC.scala 117:33]
  wire [31:0] x_13 = $signed(x_12) - $signed(_x_13_T); // @[CORDIC.scala 117:22]
  wire [19:0] _GEN_23 = fxxterm_12[31:12]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_13_T = {{12{_GEN_23[19]}},_GEN_23}; // @[CORDIC.scala 118:26]
  wire [31:0] y_13 = $signed(_y_13_T) + $signed(y_12); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_52 = $signed(theta_13) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_55 = 32'sh0 - $signed(x_13); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_13 = $signed(theta_13) > $signed(io_in_z0) ? $signed(_fxxterm_T_55) : $signed(x_13); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_55 = 32'sh0 - $signed(y_13); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_13 = _fxxterm_T_52 ? $signed(_fxyterm_T_55) : $signed(y_13); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_41 = 32'h0 - 32'h8000; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_14_T = _fxxterm_T_52 ? _fxthetaterm_T_41 : 32'h8000; // @[CORDIC.scala 116:44]
  wire [31:0] theta_14 = $signed(theta_13) + $signed(_theta_14_T); // @[CORDIC.scala 116:30]
  wire [18:0] _GEN_24 = fxyterm_13[31:13]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_14_T = {{13{_GEN_24[18]}},_GEN_24}; // @[CORDIC.scala 117:33]
  wire [31:0] x_14 = $signed(x_13) - $signed(_x_14_T); // @[CORDIC.scala 117:22]
  wire [18:0] _GEN_25 = fxxterm_13[31:13]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_14_T = {{13{_GEN_25[18]}},_GEN_25}; // @[CORDIC.scala 118:26]
  wire [31:0] y_14 = $signed(_y_14_T) + $signed(y_13); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_56 = $signed(theta_14) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_59 = 32'sh0 - $signed(x_14); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_14 = $signed(theta_14) > $signed(io_in_z0) ? $signed(_fxxterm_T_59) : $signed(x_14); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_59 = 32'sh0 - $signed(y_14); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_14 = _fxxterm_T_56 ? $signed(_fxyterm_T_59) : $signed(y_14); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_44 = 32'h0 - 32'h4000; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_15_T = _fxxterm_T_56 ? _fxthetaterm_T_44 : 32'h4000; // @[CORDIC.scala 116:44]
  wire [31:0] theta_15 = $signed(theta_14) + $signed(_theta_15_T); // @[CORDIC.scala 116:30]
  wire [17:0] _GEN_26 = fxyterm_14[31:14]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_15_T = {{14{_GEN_26[17]}},_GEN_26}; // @[CORDIC.scala 117:33]
  wire [31:0] x_15 = $signed(x_14) - $signed(_x_15_T); // @[CORDIC.scala 117:22]
  wire [17:0] _GEN_27 = fxxterm_14[31:14]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_15_T = {{14{_GEN_27[17]}},_GEN_27}; // @[CORDIC.scala 118:26]
  wire [31:0] y_15 = $signed(_y_15_T) + $signed(y_14); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_60 = $signed(theta_15) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_63 = 32'sh0 - $signed(x_15); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_15 = $signed(theta_15) > $signed(io_in_z0) ? $signed(_fxxterm_T_63) : $signed(x_15); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_63 = 32'sh0 - $signed(y_15); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_15 = _fxxterm_T_60 ? $signed(_fxyterm_T_63) : $signed(y_15); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_47 = 32'h0 - 32'h2000; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_16_T = _fxxterm_T_60 ? _fxthetaterm_T_47 : 32'h2000; // @[CORDIC.scala 116:44]
  wire [31:0] theta_16 = $signed(theta_15) + $signed(_theta_16_T); // @[CORDIC.scala 116:30]
  wire [16:0] _GEN_28 = fxyterm_15[31:15]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_16_T = {{15{_GEN_28[16]}},_GEN_28}; // @[CORDIC.scala 117:33]
  wire [31:0] x_16 = $signed(x_15) - $signed(_x_16_T); // @[CORDIC.scala 117:22]
  wire [16:0] _GEN_29 = fxxterm_15[31:15]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_16_T = {{15{_GEN_29[16]}},_GEN_29}; // @[CORDIC.scala 118:26]
  wire [31:0] y_16 = $signed(_y_16_T) + $signed(y_15); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_64 = $signed(theta_16) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_67 = 32'sh0 - $signed(x_16); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_16 = $signed(theta_16) > $signed(io_in_z0) ? $signed(_fxxterm_T_67) : $signed(x_16); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_67 = 32'sh0 - $signed(y_16); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_16 = _fxxterm_T_64 ? $signed(_fxyterm_T_67) : $signed(y_16); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_50 = 32'h0 - 32'h1000; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_17_T = _fxxterm_T_64 ? _fxthetaterm_T_50 : 32'h1000; // @[CORDIC.scala 116:44]
  wire [31:0] theta_17 = $signed(theta_16) + $signed(_theta_17_T); // @[CORDIC.scala 116:30]
  wire [15:0] _GEN_30 = fxyterm_16[31:16]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_17_T = {{16{_GEN_30[15]}},_GEN_30}; // @[CORDIC.scala 117:33]
  wire [31:0] x_17 = $signed(x_16) - $signed(_x_17_T); // @[CORDIC.scala 117:22]
  wire [15:0] _GEN_31 = fxxterm_16[31:16]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_17_T = {{16{_GEN_31[15]}},_GEN_31}; // @[CORDIC.scala 118:26]
  wire [31:0] y_17 = $signed(_y_17_T) + $signed(y_16); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_68 = $signed(theta_17) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_71 = 32'sh0 - $signed(x_17); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_17 = $signed(theta_17) > $signed(io_in_z0) ? $signed(_fxxterm_T_71) : $signed(x_17); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_71 = 32'sh0 - $signed(y_17); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_17 = _fxxterm_T_68 ? $signed(_fxyterm_T_71) : $signed(y_17); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_53 = 32'h0 - 32'h800; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_18_T = _fxxterm_T_68 ? _fxthetaterm_T_53 : 32'h800; // @[CORDIC.scala 116:44]
  wire [31:0] theta_18 = $signed(theta_17) + $signed(_theta_18_T); // @[CORDIC.scala 116:30]
  wire [14:0] _GEN_32 = fxyterm_17[31:17]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_18_T = {{17{_GEN_32[14]}},_GEN_32}; // @[CORDIC.scala 117:33]
  wire [31:0] x_18 = $signed(x_17) - $signed(_x_18_T); // @[CORDIC.scala 117:22]
  wire [14:0] _GEN_33 = fxxterm_17[31:17]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_18_T = {{17{_GEN_33[14]}},_GEN_33}; // @[CORDIC.scala 118:26]
  wire [31:0] y_18 = $signed(_y_18_T) + $signed(y_17); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_72 = $signed(theta_18) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_75 = 32'sh0 - $signed(x_18); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_18 = $signed(theta_18) > $signed(io_in_z0) ? $signed(_fxxterm_T_75) : $signed(x_18); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_75 = 32'sh0 - $signed(y_18); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_18 = _fxxterm_T_72 ? $signed(_fxyterm_T_75) : $signed(y_18); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_56 = 32'h0 - 32'h400; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_19_T = _fxxterm_T_72 ? _fxthetaterm_T_56 : 32'h400; // @[CORDIC.scala 116:44]
  wire [31:0] theta_19 = $signed(theta_18) + $signed(_theta_19_T); // @[CORDIC.scala 116:30]
  wire [13:0] _GEN_34 = fxyterm_18[31:18]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_19_T = {{18{_GEN_34[13]}},_GEN_34}; // @[CORDIC.scala 117:33]
  wire [31:0] x_19 = $signed(x_18) - $signed(_x_19_T); // @[CORDIC.scala 117:22]
  wire [13:0] _GEN_35 = fxxterm_18[31:18]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_19_T = {{18{_GEN_35[13]}},_GEN_35}; // @[CORDIC.scala 118:26]
  wire [31:0] y_19 = $signed(_y_19_T) + $signed(y_18); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_76 = $signed(theta_19) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_79 = 32'sh0 - $signed(x_19); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_19 = $signed(theta_19) > $signed(io_in_z0) ? $signed(_fxxterm_T_79) : $signed(x_19); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_79 = 32'sh0 - $signed(y_19); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_19 = _fxxterm_T_76 ? $signed(_fxyterm_T_79) : $signed(y_19); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_59 = 32'h0 - 32'h200; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_20_T = _fxxterm_T_76 ? _fxthetaterm_T_59 : 32'h200; // @[CORDIC.scala 116:44]
  wire [31:0] theta_20 = $signed(theta_19) + $signed(_theta_20_T); // @[CORDIC.scala 116:30]
  wire [12:0] _GEN_36 = fxyterm_19[31:19]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_20_T = {{19{_GEN_36[12]}},_GEN_36}; // @[CORDIC.scala 117:33]
  wire [31:0] x_20 = $signed(x_19) - $signed(_x_20_T); // @[CORDIC.scala 117:22]
  wire [12:0] _GEN_37 = fxxterm_19[31:19]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_20_T = {{19{_GEN_37[12]}},_GEN_37}; // @[CORDIC.scala 118:26]
  wire [31:0] y_20 = $signed(_y_20_T) + $signed(y_19); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_80 = $signed(theta_20) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_83 = 32'sh0 - $signed(x_20); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_20 = $signed(theta_20) > $signed(io_in_z0) ? $signed(_fxxterm_T_83) : $signed(x_20); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_83 = 32'sh0 - $signed(y_20); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_20 = _fxxterm_T_80 ? $signed(_fxyterm_T_83) : $signed(y_20); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_62 = 32'h0 - 32'h100; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_21_T = _fxxterm_T_80 ? _fxthetaterm_T_62 : 32'h100; // @[CORDIC.scala 116:44]
  wire [31:0] theta_21 = $signed(theta_20) + $signed(_theta_21_T); // @[CORDIC.scala 116:30]
  wire [11:0] _GEN_38 = fxyterm_20[31:20]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_21_T = {{20{_GEN_38[11]}},_GEN_38}; // @[CORDIC.scala 117:33]
  wire [31:0] x_21 = $signed(x_20) - $signed(_x_21_T); // @[CORDIC.scala 117:22]
  wire [11:0] _GEN_39 = fxxterm_20[31:20]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_21_T = {{20{_GEN_39[11]}},_GEN_39}; // @[CORDIC.scala 118:26]
  wire [31:0] y_21 = $signed(_y_21_T) + $signed(y_20); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_84 = $signed(theta_21) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_87 = 32'sh0 - $signed(x_21); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_21 = $signed(theta_21) > $signed(io_in_z0) ? $signed(_fxxterm_T_87) : $signed(x_21); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_87 = 32'sh0 - $signed(y_21); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_21 = _fxxterm_T_84 ? $signed(_fxyterm_T_87) : $signed(y_21); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_65 = 32'h0 - 32'h80; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_22_T = _fxxterm_T_84 ? _fxthetaterm_T_65 : 32'h80; // @[CORDIC.scala 116:44]
  wire [31:0] theta_22 = $signed(theta_21) + $signed(_theta_22_T); // @[CORDIC.scala 116:30]
  wire [10:0] _GEN_40 = fxyterm_21[31:21]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_22_T = {{21{_GEN_40[10]}},_GEN_40}; // @[CORDIC.scala 117:33]
  wire [31:0] x_22 = $signed(x_21) - $signed(_x_22_T); // @[CORDIC.scala 117:22]
  wire [10:0] _GEN_41 = fxxterm_21[31:21]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_22_T = {{21{_GEN_41[10]}},_GEN_41}; // @[CORDIC.scala 118:26]
  wire [31:0] y_22 = $signed(_y_22_T) + $signed(y_21); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_88 = $signed(theta_22) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_91 = 32'sh0 - $signed(x_22); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_22 = $signed(theta_22) > $signed(io_in_z0) ? $signed(_fxxterm_T_91) : $signed(x_22); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_91 = 32'sh0 - $signed(y_22); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_22 = _fxxterm_T_88 ? $signed(_fxyterm_T_91) : $signed(y_22); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_68 = 32'h0 - 32'h40; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_23_T = _fxxterm_T_88 ? _fxthetaterm_T_68 : 32'h40; // @[CORDIC.scala 116:44]
  wire [31:0] theta_23 = $signed(theta_22) + $signed(_theta_23_T); // @[CORDIC.scala 116:30]
  wire [9:0] _GEN_42 = fxyterm_22[31:22]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_23_T = {{22{_GEN_42[9]}},_GEN_42}; // @[CORDIC.scala 117:33]
  wire [31:0] x_23 = $signed(x_22) - $signed(_x_23_T); // @[CORDIC.scala 117:22]
  wire [9:0] _GEN_43 = fxxterm_22[31:22]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_23_T = {{22{_GEN_43[9]}},_GEN_43}; // @[CORDIC.scala 118:26]
  wire [31:0] y_23 = $signed(_y_23_T) + $signed(y_22); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_92 = $signed(theta_23) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_95 = 32'sh0 - $signed(x_23); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_23 = $signed(theta_23) > $signed(io_in_z0) ? $signed(_fxxterm_T_95) : $signed(x_23); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_95 = 32'sh0 - $signed(y_23); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_23 = _fxxterm_T_92 ? $signed(_fxyterm_T_95) : $signed(y_23); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_71 = 32'h0 - 32'h20; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_24_T = _fxxterm_T_92 ? _fxthetaterm_T_71 : 32'h20; // @[CORDIC.scala 116:44]
  wire [31:0] theta_24 = $signed(theta_23) + $signed(_theta_24_T); // @[CORDIC.scala 116:30]
  wire [8:0] _GEN_44 = fxyterm_23[31:23]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_24_T = {{23{_GEN_44[8]}},_GEN_44}; // @[CORDIC.scala 117:33]
  wire [31:0] x_24 = $signed(x_23) - $signed(_x_24_T); // @[CORDIC.scala 117:22]
  wire [8:0] _GEN_45 = fxxterm_23[31:23]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_24_T = {{23{_GEN_45[8]}},_GEN_45}; // @[CORDIC.scala 118:26]
  wire [31:0] y_24 = $signed(_y_24_T) + $signed(y_23); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_96 = $signed(theta_24) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_99 = 32'sh0 - $signed(x_24); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_24 = $signed(theta_24) > $signed(io_in_z0) ? $signed(_fxxterm_T_99) : $signed(x_24); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_99 = 32'sh0 - $signed(y_24); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_24 = _fxxterm_T_96 ? $signed(_fxyterm_T_99) : $signed(y_24); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_74 = 32'h0 - 32'h10; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_25_T = _fxxterm_T_96 ? _fxthetaterm_T_74 : 32'h10; // @[CORDIC.scala 116:44]
  wire [31:0] theta_25 = $signed(theta_24) + $signed(_theta_25_T); // @[CORDIC.scala 116:30]
  wire [7:0] _GEN_46 = fxyterm_24[31:24]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_25_T = {{24{_GEN_46[7]}},_GEN_46}; // @[CORDIC.scala 117:33]
  wire [31:0] x_25 = $signed(x_24) - $signed(_x_25_T); // @[CORDIC.scala 117:22]
  wire [7:0] _GEN_47 = fxxterm_24[31:24]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_25_T = {{24{_GEN_47[7]}},_GEN_47}; // @[CORDIC.scala 118:26]
  wire [31:0] y_25 = $signed(_y_25_T) + $signed(y_24); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_100 = $signed(theta_25) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_103 = 32'sh0 - $signed(x_25); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_25 = $signed(theta_25) > $signed(io_in_z0) ? $signed(_fxxterm_T_103) : $signed(x_25); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_103 = 32'sh0 - $signed(y_25); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_25 = _fxxterm_T_100 ? $signed(_fxyterm_T_103) : $signed(y_25); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_77 = 32'h0 - 32'h8; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_26_T = _fxxterm_T_100 ? _fxthetaterm_T_77 : 32'h8; // @[CORDIC.scala 116:44]
  wire [31:0] theta_26 = $signed(theta_25) + $signed(_theta_26_T); // @[CORDIC.scala 116:30]
  wire [6:0] _GEN_48 = fxyterm_25[31:25]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_26_T = {{25{_GEN_48[6]}},_GEN_48}; // @[CORDIC.scala 117:33]
  wire [31:0] x_26 = $signed(x_25) - $signed(_x_26_T); // @[CORDIC.scala 117:22]
  wire [6:0] _GEN_49 = fxxterm_25[31:25]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_26_T = {{25{_GEN_49[6]}},_GEN_49}; // @[CORDIC.scala 118:26]
  wire [31:0] y_26 = $signed(_y_26_T) + $signed(y_25); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_104 = $signed(theta_26) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_107 = 32'sh0 - $signed(x_26); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_26 = $signed(theta_26) > $signed(io_in_z0) ? $signed(_fxxterm_T_107) : $signed(x_26); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_107 = 32'sh0 - $signed(y_26); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_26 = _fxxterm_T_104 ? $signed(_fxyterm_T_107) : $signed(y_26); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_80 = 32'h0 - 32'h4; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_27_T = _fxxterm_T_104 ? _fxthetaterm_T_80 : 32'h4; // @[CORDIC.scala 116:44]
  wire [31:0] theta_27 = $signed(theta_26) + $signed(_theta_27_T); // @[CORDIC.scala 116:30]
  wire [5:0] _GEN_50 = fxyterm_26[31:26]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_27_T = {{26{_GEN_50[5]}},_GEN_50}; // @[CORDIC.scala 117:33]
  wire [31:0] x_27 = $signed(x_26) - $signed(_x_27_T); // @[CORDIC.scala 117:22]
  wire [5:0] _GEN_51 = fxxterm_26[31:26]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_27_T = {{26{_GEN_51[5]}},_GEN_51}; // @[CORDIC.scala 118:26]
  wire [31:0] y_27 = $signed(_y_27_T) + $signed(y_26); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_108 = $signed(theta_27) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_111 = 32'sh0 - $signed(x_27); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_27 = $signed(theta_27) > $signed(io_in_z0) ? $signed(_fxxterm_T_111) : $signed(x_27); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_111 = 32'sh0 - $signed(y_27); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_27 = _fxxterm_T_108 ? $signed(_fxyterm_T_111) : $signed(y_27); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_83 = 32'h0 - 32'h2; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_28_T = _fxxterm_T_108 ? _fxthetaterm_T_83 : 32'h2; // @[CORDIC.scala 116:44]
  wire [31:0] theta_28 = $signed(theta_27) + $signed(_theta_28_T); // @[CORDIC.scala 116:30]
  wire [4:0] _GEN_52 = fxyterm_27[31:27]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_28_T = {{27{_GEN_52[4]}},_GEN_52}; // @[CORDIC.scala 117:33]
  wire [31:0] x_28 = $signed(x_27) - $signed(_x_28_T); // @[CORDIC.scala 117:22]
  wire [4:0] _GEN_53 = fxxterm_27[31:27]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_28_T = {{27{_GEN_53[4]}},_GEN_53}; // @[CORDIC.scala 118:26]
  wire [31:0] y_28 = $signed(_y_28_T) + $signed(y_27); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_112 = $signed(theta_28) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_115 = 32'sh0 - $signed(x_28); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_28 = $signed(theta_28) > $signed(io_in_z0) ? $signed(_fxxterm_T_115) : $signed(x_28); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_115 = 32'sh0 - $signed(y_28); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_28 = _fxxterm_T_112 ? $signed(_fxyterm_T_115) : $signed(y_28); // @[CORDIC.scala 113:22]
  wire [31:0] _fxthetaterm_T_86 = 32'h0 - 32'h1; // @[CORDIC.scala 114:46]
  wire [31:0] _theta_29_T = _fxxterm_T_112 ? _fxthetaterm_T_86 : 32'h1; // @[CORDIC.scala 116:44]
  wire [31:0] theta_29 = $signed(theta_28) + $signed(_theta_29_T); // @[CORDIC.scala 116:30]
  wire [3:0] _GEN_54 = fxyterm_28[31:28]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_29_T = {{28{_GEN_54[3]}},_GEN_54}; // @[CORDIC.scala 117:33]
  wire [31:0] x_29 = $signed(x_28) - $signed(_x_29_T); // @[CORDIC.scala 117:22]
  wire [3:0] _GEN_55 = fxxterm_28[31:28]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_29_T = {{28{_GEN_55[3]}},_GEN_55}; // @[CORDIC.scala 118:26]
  wire [31:0] y_29 = $signed(_y_29_T) + $signed(y_28); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_116 = $signed(theta_29) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_119 = 32'sh0 - $signed(x_29); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_29 = $signed(theta_29) > $signed(io_in_z0) ? $signed(_fxxterm_T_119) : $signed(x_29); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_119 = 32'sh0 - $signed(y_29); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_29 = _fxxterm_T_116 ? $signed(_fxyterm_T_119) : $signed(y_29); // @[CORDIC.scala 113:22]
  wire [32:0] _theta_30_T_1 = {{1{theta_29[31]}},theta_29}; // @[CORDIC.scala 116:30]
  wire [31:0] theta_30 = _theta_30_T_1[31:0]; // @[CORDIC.scala 116:30]
  wire [2:0] _GEN_56 = fxyterm_29[31:29]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_30_T = {{29{_GEN_56[2]}},_GEN_56}; // @[CORDIC.scala 117:33]
  wire [31:0] x_30 = $signed(x_29) - $signed(_x_30_T); // @[CORDIC.scala 117:22]
  wire [2:0] _GEN_57 = fxxterm_29[31:29]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_30_T = {{29{_GEN_57[2]}},_GEN_57}; // @[CORDIC.scala 118:26]
  wire [31:0] y_30 = $signed(_y_30_T) + $signed(y_29); // @[CORDIC.scala 118:46]
  wire  _fxxterm_T_120 = $signed(theta_30) > $signed(io_in_z0); // @[CORDIC.scala 112:32]
  wire [31:0] _fxxterm_T_123 = 32'sh0 - $signed(x_30); // @[CORDIC.scala 112:42]
  wire [31:0] fxxterm_30 = $signed(theta_30) > $signed(io_in_z0) ? $signed(_fxxterm_T_123) : $signed(x_30); // @[CORDIC.scala 112:22]
  wire [31:0] _fxyterm_T_123 = 32'sh0 - $signed(y_30); // @[CORDIC.scala 113:42]
  wire [31:0] fxyterm_30 = _fxxterm_T_120 ? $signed(_fxyterm_T_123) : $signed(y_30); // @[CORDIC.scala 113:22]
  wire [1:0] _GEN_58 = fxyterm_30[31:30]; // @[CORDIC.scala 117:33]
  wire [31:0] _x_31_T = {{30{_GEN_58[1]}},_GEN_58}; // @[CORDIC.scala 117:33]
  wire [1:0] _GEN_59 = fxxterm_30[31:30]; // @[CORDIC.scala 118:26]
  wire [31:0] _y_31_T = {{30{_GEN_59[1]}},_GEN_59}; // @[CORDIC.scala 118:26]
  FloatToFixed32 tofixedx0 ( // @[CORDIC.scala 63:25]
    .io_in(tofixedx0_io_in),
    .io_out(tofixedx0_io_out)
  );
  FloatToFixed32 tofixedy0 ( // @[CORDIC.scala 64:25]
    .io_in(tofixedy0_io_in),
    .io_out(tofixedy0_io_out)
  );
  FixedToFloat32 tofloatxout ( // @[CORDIC.scala 123:27]
    .io_in(tofloatxout_io_in),
    .io_out(tofloatxout_io_out)
  );
  FixedToFloat32 tofloatyout ( // @[CORDIC.scala 124:27]
    .io_in(tofloatyout_io_in),
    .io_out(tofloatyout_io_out)
  );
  FixedToFloat32 tofloatzout ( // @[CORDIC.scala 125:27]
    .io_in(tofloatzout_io_in),
    .io_out(tofloatzout_io_out)
  );
  assign io_out_x = tofloatxout_io_out; // @[CORDIC.scala 132:12]
  assign io_out_mode = io_in_mode[1:0]; // @[CORDIC.scala 108:12 74:19]
  assign tofixedx0_io_in = 32'h3f1b74ee; // @[CORDIC.scala 67:19]
  assign tofixedy0_io_in = 32'h0; // @[CORDIC.scala 68:19]
  assign tofloatxout_io_in = $signed(x_30) - $signed(_x_31_T); // @[CORDIC.scala 128:30]
  assign tofloatyout_io_in = $signed(_y_31_T) + $signed(y_30); // @[CORDIC.scala 129:30]
  assign tofloatzout_io_in = io_in_z0; // @[CORDIC.scala 130:32]
endmodule
module Sin(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out
);
  wire [31:0] tofixedz0_io_in; // @[Sin.scala 23:25]
  wire [31:0] tofixedz0_io_out; // @[Sin.scala 23:25]
  wire [31:0] cordic_io_in_z0; // @[Sin.scala 27:22]
  wire [31:0] cordic_io_in_mode; // @[Sin.scala 27:22]
  wire [31:0] cordic_io_out_x; // @[Sin.scala 27:22]
  wire [1:0] cordic_io_out_mode; // @[Sin.scala 27:22]
  wire [31:0] adjangle = 32'sh1921fb60 - $signed(tofixedz0_io_out); // @[Sin.scala 43:29]
  wire [31:0] _theta_T_3 = $signed(adjangle) + 32'sh6487ed80; // @[Sin.scala 44:44]
  wire [31:0] theta = $signed(adjangle) < 32'sh0 ? $signed(_theta_T_3) : $signed(adjangle); // @[Sin.scala 44:18]
  wire  _T_3 = $signed(theta) > 32'sh1921fb60 & $signed(theta) < 32'sh4b65f200; // @[Sin.scala 50:33]
  wire [1:0] _GEN_1 = $signed(theta) > 32'sh4b65f200 ? 2'h2 : {{1'd0}, _T_3}; // @[Sin.scala 48:33 49:23]
  wire [31:0] _cordic_io_in_z0_T_3 = $signed(theta) - 32'sh6487ed80; // @[Sin.scala 58:41]
  wire [31:0] _cordic_io_in_z0_T_7 = 32'sh3243f6c0 - $signed(theta); // @[Sin.scala 61:37]
  wire  _io_out_T_1 = ~cordic_io_out_x[31]; // @[Sin.scala 62:15]
  wire [31:0] _io_out_T_3 = {_io_out_T_1,cordic_io_out_x[30:0]}; // @[Sin.scala 62:36]
  wire [31:0] _cordic_io_in_z0_T_8 = $signed(adjangle) < 32'sh0 ? $signed(_theta_T_3) : $signed(adjangle); // @[Sin.scala 65:30]
  wire [31:0] _GEN_2 = cordic_io_out_mode == 2'h1 ? _cordic_io_in_z0_T_7 : _cordic_io_in_z0_T_8; // @[Sin.scala 60:30 61:21 65:21]
  wire [31:0] _GEN_3 = cordic_io_out_mode == 2'h1 ? _io_out_T_3 : cordic_io_out_x; // @[Sin.scala 60:30 62:12 66:12]
  FloatToFixed32 tofixedz0 ( // @[Sin.scala 23:25]
    .io_in(tofixedz0_io_in),
    .io_out(tofixedz0_io_out)
  );
  CORDIC cordic ( // @[Sin.scala 27:22]
    .io_in_z0(cordic_io_in_z0),
    .io_in_mode(cordic_io_in_mode),
    .io_out_x(cordic_io_out_x),
    .io_out_mode(cordic_io_out_mode)
  );
  assign io_out = cordic_io_out_mode == 2'h2 ? cordic_io_out_x : _GEN_3; // @[Sin.scala 57:24 59:12]
  assign tofixedz0_io_in = io_in; // @[Sin.scala 24:19]
  assign cordic_io_in_z0 = cordic_io_out_mode == 2'h2 ? _cordic_io_in_z0_T_3 : _GEN_2; // @[Sin.scala 57:24 58:21]
  assign cordic_io_in_mode = {{30'd0}, _GEN_1};
endmodule

